.include "./bin_0_nch_modified.lib"

.option verbose=1

* IV VDS Simulation netlist for NMOS using MODIFIED model
* Model: sky130_fd_pr__nfet_01v8__model.0
.param nf=1
.param w=1.26
.param l=0.15

M1 net1 VGS GND GND sky130_fd_pr__nfet_01v8__model.0 L=0.15 W=1.26 nf=1 ad='int((nf+1)/2)*w/nf*0.29' as='int((nf+2)/2)*w/nf*0.29'
+pd='2*int((nf+1)/2)*(w/nf+0.29)' ps='2*int((nf+2)/2)*(w/nf+0.29)' nrd='0.29/w' nrs='0.29/w' sa=0 sb=0 sd=0
VGATE VGS GND 0
VDRAIN VDS GND 0
vdsM VDS net1 0

.save i(vdsm)

.control
save all
let vgsval = 0
let step = 0.6
while vgsval <= 1.8
    echo Sweeping VGS = $&vgsval
    alter VGATE = $&vgsval
    dc VDRAIN 0 1.8 0.1
    wrdata results_IV_ID_vs_VDS_for_VG_sweep/n_mosfet_id_vs_vsd_{$&vgsval}.csv V(VDS) I(VDRAIN) I(VDSM)
    let vgsval = $&vgsval + $&step
end
write results_IV_ID_vs_VDS_for_VG_sweep/IV_IDS_vs_VDS.raw
.endc

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/designs/sky130A/libs.tech/ngspice/corners/tt/spice
.include /foss/designs/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/designs/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/designs/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

.GLOBAL GND
.end
