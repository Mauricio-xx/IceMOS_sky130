.include "./bin_0_nch_modified.lib"

.option verbose=1

* IV VDS Simulation netlist for device nch using MODIFIED model
* Model: sky130_fd_pr__nfet_01v8__model.0
* Parameter definitions for device dimensions
.param nf=1
.param w=1
.param l=0.15

* MOSFET instance using the defined parameters
M1 net1 VGS GND GND sky130_fd_pr__nfet_01v8__model.0 L=1 W=1 nf=1 ad='int((nf+1)/2)*W/nf*0.29' as='int((nf+2)/2)*W/nf*0.29' pd='2*int((nf+1)/2)*(W/nf+0.29)' 
+ ps='2*int((nf+2)/2)*(W/nf+0.29)' nrd='0.29/W' nrs='0.29/W' sa=0 sb=0 sd=0 m=1

VGATE VGS GND 0
VDRAIN VDS GND 0
vdsM VDS net1 0

.save i(vdsm)

.control
save all
* op
  * Initialize VGS and step
let vgsval = 0
let step = 0.6

* Sweep VGS from 0V to 1.8V in steps of 0.6V
while vgsval <= 1.8
    echo Sweeping VGS = $&vgsval
    alter VGATE = $&vgsval
    dc VDRAIN 0 1.8 0.1
    wrdata sweep_IV_results/mosfet_vds_vs_id_{$&vgsval}.csv V(VDS) I(VDRAIN) I(VDSM)
    let vgsval = $&vgsval + $&step
end
write IV_IDS_vs_VDS.raw
.endc

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

.GLOBAL GND
.end
