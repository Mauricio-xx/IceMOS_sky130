** sch_path: /foss/designs/IceMOS_sky130/circuits/copys_to_develop_pmos/IV_ISD_vs_VSD?.sch
**.subckt IV_ISD_vs_VSD?
VGATE VGS GND 0
VSOURCE VSD GND 0
vsdM VSD net1 0
.save i(vsdm)
XM2 GND VGS net1 GND sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code



*.control
*save all
*op
    * VDS sweep and VGS sweep
*    dc VDRAIN 0 1.8 0.01 VGATE 0 1.8 0.6
    * Save the results
*    wrdata mosfet_vds_vs_is.csv V(VGS) I(VDRAIN)
*.endc



.control
save all
op
  * Barrido de VGS de 0V a 1.8V en pasos de 0.6V
  foreach vgs 0 0.1 0.2 0.3 0.4 0.5 0.6 1.2 1.8
    * Cambiar VGS a $vgs
    alter VGATE dc=$vgs
    * Barrido de VSD de 0V a 1.8V en pasos de 0.1V
    dc VSOURCE 0 1.8 0.1
    * Guardar los resultados en un archivo
    wrdata mosfet_vsd_vs_is_{$vgs}.csv V(VGS) I(VSOURCE) I(vsdM)

  end
write IV_ISD_vs_VSD.raw
.endc



.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends
.GLOBAL GND
.end
