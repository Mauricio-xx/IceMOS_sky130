.include "./bin_40_nch_original.lib"

.option verbose=1

*set temperature for simulation
*if this file is 'ORIGINAL' temp is set to 27C
*if this file is 'MODIFIED' temp is -269C (4K)
.temp 27

* IV VDS Simulation netlist for NMOS using ORIGINAL model
* Model: sky130_fd_pr__nfet_01v8__model.40
.param nf=1
.param w=0.42
.param l=0.15

M1 net1 VGS GND GND sky130_fd_pr__nfet_01v8__model.40 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2)*w/nf*0.29' as='int((nf+2)/2)*w/nf*0.29'
+pd='2*int((nf+1)/2)*(w/nf+0.29)' ps='2*int((nf+2)/2)*(w/nf+0.29)' nrd='0.29/w' nrs='0.29/w' sa=0 sb=0 sd=0
VGATE VGS GND 0
VDRAIN VDS GND 0
vdsM VDS net1 0

.save i(vdsm)

.control
save all
let vgsval = 0.9
let step = 0.3
while vgsval <= 1.8
    echo Sweeping VGS = $&vgsval
    alter VGATE = $&vgsval
    dc VDRAIN 0.0 1.8 0.1
    wrdata results_IV_IDS_vs_VDS_for_VG_sweep/n_mosfet_id_vs_vsd_{$&vgsval}.csv V(VDS) I(VDRAIN) I(VDSM)
    write results_IV_IDS_vs_VDS_for_VG_sweep/n_mosfet_id_vs_vsd_{$&vgsval}.raw
    let vgsval = $&vgsval + $&step
end

.endc


.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice
.GLOBAL GND
.end
