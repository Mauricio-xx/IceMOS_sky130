** sch_path: /foss/designs/Endurance_Cryo_ToolBox/src/exp/sky130/nch/IV_current_vs_vdrain/IV_IDS_vs_VDS.sch
**.subckt IV_IDS_vs_VDS
XM1 net1 VGS GND GND sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
VGATE VGS GND 0
VDRAIN VDS GND 0
vdsM VDS net1 0
.save i(vdsm)
**** begin user architecture code



.control
save all
* op
  * Initialize VGS and step
let vgsval = 0
let step = 0.6

* Sweep VGS from 0V to 1.8V in steps of 0.6V
while vgsval <= 1.8

	echo Sweeping VGS = $&vgsval

	* pass vgs to VGATE (circuit level)
	alter VGATE = $&vgsval
	* Sweep VDS from 0V to 1.8V in steps of 0.1V
    	dc VDRAIN 0 1.8 0.1

    	* Save the results to a file
    	wrdata mosfet_vds_vs_id_{$&vgsval}.csv V(VDS) I(VDRAIN) I(VDSM)

    	* Increment VGS
    	let vgsval = $&vgsval + $&step
end

write IV_IDS_vs_VDS.raw
.endc




.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
