** sch_path: /foss/designs/Endurance_Cryo_ToolBox/src/exp/sky130/nch/IV_nmos.sch
**.subckt IV_nmos
VGATE net1 GND 0
XM1 net2 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V1 V1 GND 1.8
V1_meas V1 net2 0
.save i(v1_meas)
**** begin user architecture code

.control
save all
*op
*write  IV_nmos.raw

* Perform DC sweep for V1 from 0V to 1.8V in steps of 0.1V
dc VGATE 0 1.8 0.1

*print I(v1)

write IV_nmos.raw
wrdata IV_nmos.csv I(v1)


.endc



.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
