.include "./bin_40_nch_modified.lib"

.option verbose=1

*set temperature for simulation
*if this file is 'ORIGINAL' temp is set to 27C
*if this file is 'MODIFIED' temp is -269C (4K)
.temp -269

* IV Simulation netlist for device nch using MODIFIED model
* Model: sky130_fd_pr__nfet_01v8__model.40
.param nf=1
.param w=0.42
.param l=0.15

VGATE_src net1 GND 0
M1 net2 net1 0 0 sky130_fd_pr__nfet_01v8__model.40 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2)*W/nf*0.29' as='int((nf+2)/2)*W/nf*0.29'
+pd='2*int((nf+1)/2)*(W/nf+0.29)' ps='2*int((nf+2)/2)*(W/nf+0.29)' nrd='0.29/W' nrs='0.29/W' sa=0 sb=0 sd=0
V1 V1 GND 1.8
V1_meas V1 net2 0
.save i(V1_meas)

.control
  save all
  dc VGATE_src 0.0 1.8 0.01
  write results_IV_ID_vs_VG/IV_ID_vs_VG.raw
  wrdata results_IV_ID_vs_VG/IV_ID_vs_VG.csv I(V1_meas)
  *showmod M1
.endc

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

.GLOBAL GND
.end
